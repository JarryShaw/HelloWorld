// File: Verilog.v

module Verilog ();

    initial begin
        $display("Across the Great Wall, we can reach every corner in the world.")
    end

endmodule // Verilog
